* D:\Prakalp\SFAL_tool\Inv_A\Inv_A.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 1/30/2022 6:30:09 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad1_ /Vout GND GND mosfet_n		
U1  /Vdd PORT		
U3  /Vout PORT		
M3  Net-_M3-Pad1_ Net-_M1-Pad1_ /Vdd /Vdd mosfet_p		
M4  Net-_M3-Pad1_ Net-_M1-Pad1_ GND GND mosfet_n		
M5  Net-_M5-Pad1_ Net-_M3-Pad1_ /Vdd /Vdd mosfet_p		
M6  Net-_M5-Pad1_ Net-_M3-Pad1_ GND GND mosfet_n		
M7  Net-_M10-Pad2_ Net-_M5-Pad1_ /Vdd /Vdd mosfet_p		
M8  Net-_M10-Pad2_ Net-_M5-Pad1_ GND GND mosfet_n		
M9  Net-_M10-Pad1_ Net-_M10-Pad2_ /Vdd /Vdd mosfet_p		
M10  Net-_M10-Pad1_ Net-_M10-Pad2_ GND GND mosfet_n		
M11  Net-_M11-Pad1_ Net-_M10-Pad1_ /Vdd /Vdd mosfet_p		
M12  Net-_M11-Pad1_ Net-_M10-Pad1_ GND GND mosfet_n		
M13  Net-_M13-Pad1_ Net-_M11-Pad1_ /Vdd /Vdd mosfet_p		
M14  Net-_M13-Pad1_ Net-_M11-Pad1_ GND GND mosfet_n		
M15  Net-_M15-Pad1_ Net-_M13-Pad1_ /Vdd /Vdd mosfet_p		
M16  Net-_M15-Pad1_ Net-_M13-Pad1_ GND GND mosfet_n		
M17  /Vout Net-_M15-Pad1_ /Vdd /Vdd mosfet_p		
M18  /Vout Net-_M15-Pad1_ GND GND mosfet_n		
M1  Net-_M1-Pad1_ /Vout /Vdd /Vdd mosfet_p		

.end
